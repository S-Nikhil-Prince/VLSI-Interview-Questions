1)5:1 mux using 2:1 mux
2)2:1 mux using 4:1 mux
3)all 2 input logic gates(AND,OR,NAND,NOR,EX-OR,EX-NOR) using mux
4)all 3 input logic gates(AND,OR,NAND,NOR,EX-OR,EX-NOR) using mux
5)Design full adder using i) 4:1 Mux and 1 not gate   ii) 2:1 Mux only   iii) 8:1 Mux     iv) 16:1 mux
6)design 10:1 mux using 3x(4:1 Mux)
7)design 4:1 mux using decoder and trisate buffer
8)implement nand using nor and vice versa
9)implement 3:1 mux using 2:1 mux with following selection requirments 
    i)ab=00 then i0
    ii)ab=01 then i3
    iii)ab=10 then i2
10) design 2:1 mux nor gate only and also using nand gate only
11)f(a,b,c,d) = E
12)
13)